// Troy Kaufman
// tkaufman@g.hmc.edu
// 10/27/24
// This module adds the current state with a round key produced by key_expansion's key schedule

module add_round_key(input logic [127:0] state, round_key,
                     output logic [127:0] new_state);

    assign new_state = state ^ key;

endmodule

