// Troy Kaufman
// tkaufman@g.hmc.edu
// 10/27/24
// This module rotates a four byte sequence

module rot_Word(input logic [7:0] b0, b1, b2, b3,
                output logic [31:0] row_of_bytes);

    assign row_of_bytes = {b1, b2, b3, b0};

endmodule